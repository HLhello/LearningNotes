module led_ipcnt(
	clk,
	rst,
	led
);

input clk;
input rst;

output reg led;




endmodule  