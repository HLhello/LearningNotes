module speed_setting(
	clk,
	rst,
	
);

input clk;
input rst;


endmodule 