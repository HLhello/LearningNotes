module key_board(
	clk,
	rst,
	key_row,
	key_flag,
	key_value,
	key_col
);

input clk;
input rst
input [3:0]key_row;
output key_flag;
output [3:0]key_value;
output [3:0]key_col;




endmodule

