module testtteets();


endmodule 