module uart_tx(
	clk,
	rst,
	
);

input clk;
input rst;


endmodule 