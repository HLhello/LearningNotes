module key_filter(

);

endmodule

