module pwm_gen(
	clk,
	rst,
	cnt_en,
	cnt_arr,
	cnt_ccr,
	o_pwm
);

input clk;
input rst;
input cnt_en;
input [31:0]cnt_arr;
input [31:0]cnt_ccr;
output o_pwm;


endmodule 
