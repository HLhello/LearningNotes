module key_filter(
	clk,
	rst,
	key_in,
	key_flag,
	key_state
);

input clk,
input rst,
input key_in,
output reg key_flag,
output reg key_state




endmodule 
