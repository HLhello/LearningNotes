module rx_bps_gen(
	clk,
	rst,
	baud_set,
	rx_done,
	byte_en,
	sample_clk
);

input clk;
input rst;
input [2:0]baud_set;
input rx_done;
input byte_en;
output reg sample_clk;


endmodule 
