module uart_rx(
	clk,
	rst,
	
);

input clk;
input rst;


endmodule 