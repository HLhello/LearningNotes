module fsm_welcome(

);



endmodule 

