module fsm_keystate(

);

endmodule

