module tx_bps_gen(
	clk,
	rst,
	baud_set,
	tx_done,
	bps_en,
	bps_clk
);

input clk;
input rst;
input [2:0]baud_set;
input tx_done;
input bps_en;
output reg bps_clk;


endmodule 
